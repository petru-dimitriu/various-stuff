module inc(in, out);

input [31:0] in;
output [31:0] out;

assign out = in + 3'b100;

endmodule
